CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
550 540 30 70 10
1542 80 2644 963
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 1
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
1710 176 1823 273
77070354 0
0
6 Title:
5 Name:
0
0
0
71
7 Ground~
168 1413 1233 0 1 3
0 2
0
0 0 53344 0
0
5 GND13
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
631 0 0
2
42619.7 0
0
5 SIP5~
219 1440 1152 0 5 11
0 6 5 2 3 4
0
0 0 864 0
4 MCHP
-11 -43 17 -35
2 W3
-4 -34 10 -26
0
0
0
0
0
4 SIP5
11

0 1 2 3 4 5 1 2 3 4
5 0
0 0 0 0 1 0 0 0
1 J
9466 0 0
2
42619.7 1
0
10 Capacitor~
219 1314 1197 0 2 5
0 2 5
0
0 0 832 90
4 10uF
9 4 37 12
3 C15
11 -7 32 1
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 22
67 0 0 0 1 0 0 0
1 C
3266 0 0
2
42619.7 2
0
10 Capacitor~
219 1260 1197 0 2 5
0 2 5
0
0 0 832 90
5 0.1uF
5 4 40 12
3 C14
11 -6 32 2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 266
67 0 0 0 1 0 0 0
1 C
7693 0 0
2
42619.7 3
0
9 Inductor~
219 1080 1017 0 2 5
0 11 5
0
0 0 1856 0
5 4.7uH
-18 -17 17 -9
2 L1
-7 -27 7 -19
4 20mA
-14 -37 14 -29
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
3723 0 0
2
42619.7 4
0
10 Capacitor~
219 972 1170 0 2 5
0 2 12
0
0 0 832 90
4 10uF
-35 1 -7 9
3 C12
-32 -8 -11 0
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 250
67 0 0 0 1 0 0 0
1 C
3440 0 0
2
42619.7 5
0
7 Ground~
168 990 1215 0 1 3
0 2
0
0 0 53344 0
0
5 GND12
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6263 0 0
2
42619.7 6
0
7 Ground~
168 1233 1233 0 1 3
0 2
0
0 0 53344 0
0
5 GND11
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4900 0 0
2
42619.7 7
0
7 Ground~
168 1188 1302 0 1 3
0 2
0
0 0 53344 0
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8783 0 0
2
42619.7 8
0
7 Ground~
168 1125 1302 0 1 3
0 2
0
0 0 53344 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3221 0 0
2
42619.7 9
0
10 Capacitor~
219 1125 1287 0 2 5
0 2 14
0
0 0 832 90
4 22pF
9 0 37 8
3 C11
12 -9 33 -1
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 74075136
67 0 0 0 1 0 0 0
1 C
3215 0 0
2
42619.7 10
0
10 Capacitor~
219 1188 1287 0 2 5
0 2 13
0
0 0 832 90
3 1uF
11 0 32 8
3 C10
11 -10 32 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 250
67 0 0 0 1 0 0 0
1 C
7903 0 0
2
42619.7 11
0
8 Crystal~
219 1159 1269 0 2 5
0 14 13
0
0 0 832 0
9 10.000MHZ
-31 -18 32 -10
5 XTAL1
-18 -28 17 -20
0
0
11 %D %1 %2 %S
0
14 alias:XCRYSTAL
5 XTAL1
5

0 1 2 1 2 0
88 0 0 0 1 0 0 0
4 XTAL
7121 0 0
2
42619.7 12
0
7 Ground~
168 1296 1113 0 1 3
0 2
0
0 0 53344 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4484 0 0
2
42619.7 13
0
12 SPST Switch~
165 1295 1062 0 2 11
0 15 16
0
0 0 4704 90
0
2 S1
11 -6 25 2
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
5996 0 0
2
42619.7 14
0
10 Capacitor~
219 1296 1098 0 2 5
0 2 16
0
0 0 832 90
3 1uF
11 0 32 8
2 C9
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 74076532
67 0 0 0 1 0 0 0
1 C
7804 0 0
2
42619.7 15
0
2 +V
167 1350 963 0 1 3
0 5
0
0 0 53728 0
2 5V
-6 -20 8 -12
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5523 0 0
2
42619.7 16
0
7 Ground~
168 711 861 0 1 3
0 2
0
0 0 53344 0
0
5 GND26
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3330 0 0
2
5.89768e-315 0
0
10 Capacitor~
219 711 846 0 2 5
0 2 23
0
0 0 1856 90
5 4.7uF
9 0 44 8
3 C23
11 -10 32 -2
3 50V
11 -20 32 -12
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 74041768
67 0 0 0 1 0 0 0
1 C
3465 0 0
2
5.89768e-315 5.26354e-315
0
9 Schottky~
219 677 828 0 2 5
0 24 23
0
0 0 832 0
6 1N5817
-20 -18 22 -10
2 D4
-6 -28 8 -20
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
8396 0 0
2
5.89768e-315 5.30499e-315
0
4 LED~
171 1946 699 0 2 2
10 25 2
0
0 0 864 90
5 AMBER
-15 -21 20 -13
2 D2
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3685 0 0
2
5.89768e-315 5.32571e-315
0
4 LED~
171 1641 699 0 2 2
10 27 2
0
0 0 864 90
5 GREEN
-15 -21 20 -13
2 D1
-5 -31 9 -23
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
7849 0 0
2
5.89768e-315 5.34643e-315
0
2 +V
167 1894 682 0 1 3
0 25
0
0 0 53728 0
4 3.3V
-13 -20 15 -12
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6343 0 0
2
5.89768e-315 5.3568e-315
0
10 Polar Cap~
219 1841 737 0 2 5
0 25 2
0
0 0 832 270
5 220uF
9 3 44 11
2 C4
18 -6 32 2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7376 0 0
2
5.89768e-315 5.36716e-315
0
10 Capacitor~
219 1894 736 0 2 5
0 2 25
0
0 0 832 90
5 0.1uF
10 0 45 8
2 C5
19 -10 33 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9156 0 0
2
5.89768e-315 5.37752e-315
0
10 Capacitor~
219 1741 736 0 2 5
0 2 28
0
0 0 832 90
3 1uF
-30 0 -9 8
2 C6
-26 -9 -12 -1
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5776 0 0
2
5.89768e-315 5.38788e-315
0
7 Ground~
168 1795 772 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7207 0 0
2
5.89768e-315 5.39306e-315
0
7 Ground~
168 1741 772 0 1 3
0 2
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4459 0 0
2
5.89768e-315 5.39824e-315
0
2 +V
167 1741 682 0 1 3
0 28
0
0 0 53984 0
3 12V
-11 -22 10 -14
4 BATT
-13 -20 15 -12
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3760 0 0
2
5.89768e-315 5.40342e-315
0
11 Regulator3~
219 1795 727 0 3 7
0 28 2 25
0
0 0 4928 0
10 LD1117AV33
-35 -28 35 -20
2 U3
-7 -38 7 -30
0
0
14 %D %1 %2 %3 %S
0
0
6 TO-220
7

0 3 1 2 3 1 2 0
88 0 0 0 1 1 0 0
1 U
754 0 0
2
5.89768e-315 5.4086e-315
0
11 Regulator3~
219 1486 728 0 3 7
0 29 2 26
0
0 0 4928 0
5 78L05
-18 -28 17 -20
2 U2
-7 -38 7 -30
0
0
14 %D %1 %2 %3 %S
0
0
6 TO-220
7

0 3 1 2 3 1 2 0
88 0 0 0 1 1 0 0
1 U
9767 0 0
2
5.89768e-315 5.41378e-315
0
2 +V
167 1432 683 0 1 3
0 29
0
0 0 53984 0
3 10V
-11 -22 10 -14
4 BATT
-13 -20 15 -12
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7978 0 0
2
5.89768e-315 5.41896e-315
0
7 Ground~
168 1432 773 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3142 0 0
2
5.89768e-315 5.42414e-315
0
7 Ground~
168 1486 773 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3284 0 0
2
5.89768e-315 5.42933e-315
0
10 Capacitor~
219 1432 737 0 2 5
0 2 29
0
0 0 832 90
3 1uF
-30 0 -9 8
2 C1
-26 -9 -12 -1
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
659 0 0
2
5.89768e-315 5.43192e-315
0
10 Capacitor~
219 1585 737 0 2 5
0 2 26
0
0 0 832 90
5 0.1uF
10 0 45 8
2 C2
19 -10 33 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3800 0 0
2
5.89768e-315 5.43451e-315
0
10 Polar Cap~
219 1532 738 0 2 5
0 26 2
0
0 0 832 270
5 220uF
9 3 44 11
2 C3
18 -6 32 2
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6792 0 0
2
5.89768e-315 5.4371e-315
0
2 +V
167 1585 683 0 1 3
0 26
0
0 0 53728 0
2 5V
-6 -20 8 -12
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3701 0 0
2
5.89768e-315 5.43969e-315
0
7 Ground~
168 873 1095 0 1 3
0 2
0
0 0 53344 0
0
5 GND25
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6316 0 0
2
5.89768e-315 5.44228e-315
0
7 Ground~
168 810 1095 0 1 3
0 2
0
0 0 53344 0
0
5 GND24
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8734 0 0
2
5.89768e-315 5.44487e-315
0
10 Capacitor~
219 810 1080 0 2 5
0 2 30
0
0 0 832 90
4 22pF
7 0 35 8
3 C22
11 -10 32 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 26
67 0 0 0 1 0 0 0
1 C
7988 0 0
2
5.89768e-315 5.44746e-315
0
10 Capacitor~
219 873 1080 0 2 5
0 2 31
0
0 0 832 90
4 22pF
8 0 36 8
3 C21
11 -10 32 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 62
67 0 0 0 1 0 0 0
1 C
3217 0 0
2
5.89768e-315 5.45005e-315
0
8 Crystal~
219 844 1053 0 2 5
0 30 31
0
0 0 832 0
9 16.000MHZ
-32 -18 31 -10
5 XTAL2
-18 -28 17 -20
0
0
11 %D %1 %2 %S
0
14 alias:XCRYSTAL
5 XTAL1
5

0 1 2 1 2 0
88 0 0 0 1 0 0 0
4 XTAL
3965 0 0
2
5.89768e-315 5.45264e-315
0
7 Ground~
168 684 1023 0 1 3
0 2
0
0 0 53344 0
0
5 GND18
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8239 0 0
2
42619.7 17
0
4 LED~
171 684 1000 0 2 2
10 32 2
0
0 0 864 0
4 BLUE
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
828 0 0
2
42619.7 18
0
7 Ground~
168 864 915 0 1 3
0 2
0
0 0 53344 0
0
5 GND17
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6187 0 0
2
42619.7 19
0
10 Capacitor~
219 864 900 0 2 5
0 2 35
0
0 0 832 90
3 1uF
11 0 32 8
2 C8
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7107 0 0
2
42619.7 20
0
7 Ground~
168 747 897 0 1 3
0 2
0
0 0 53344 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6433 0 0
2
42619.7 21
0
10 Capacitor~
219 747 882 0 2 5
0 2 35
0
0 0 832 90
5 100nF
9 0 44 8
2 C7
19 -10 33 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
8559 0 0
2
42619.7 22
0
2 +V
167 801 847 0 1 3
0 35
0
0 0 53728 0
2 5V
-6 -20 8 -12
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3674 0 0
2
42619.7 23
0
7 Ground~
168 783 1023 0 1 3
0 2
0
0 0 53344 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5697 0 0
2
42619.7 24
0
5 DB-9~
219 625 864 0 9 19
0 45 46 47 48 49 33 34 2 24
0
0 0 2656 0
4 CONN
30 2 58 10
2 J1
-7 -50 7 -42
0
0
0
0
0
5 DB9/F
19

0 1 2 3 4 5 -13589035 -13589039 -195123 -8605027
1 2 3 4 5 -13589035 -13589039 -195123 -8605027 0
0 0 0 512 1 1 0 0
1 J
3805 0 0
2
42619.7 25
0
7 Ground~
168 666 918 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5219 0 0
2
42619.7 26
0
2 +V
167 711 783 0 1 3
0 23
0
0 0 54112 0
3 12V
-11 -13 10 -5
4 BATT
-14 -22 14 -14
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3795 0 0
2
42619.7 27
0
10 Capacitor~
219 1179 639 0 2 5
0 2 38
0
0 0 1856 90
3 1uF
-29 3 -8 11
3 C17
-29 -7 -8 1
3 50V
-29 14 -8 22
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 62
67 0 0 0 1 0 0 0
1 C
3637 0 0
2
5.89768e-315 5.45523e-315
0
2 +V
167 1179 585 0 1 3
0 38
0
0 0 53984 0
3 12V
-9 -19 12 -11
4 BATT
-13 -19 15 -11
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3226 0 0
2
5.89768e-315 5.45782e-315
0
10 Capacitor~
219 1308 666 0 2 5
0 2 39
0
0 0 1856 180
5 0.1uF
-18 -18 17 -10
3 C20
-11 -28 10 -20
3 20V
-10 11 11 19
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 22
67 0 0 0 1 0 0 0
1 C
6966 0 0
2
5.89768e-315 5.46041e-315
0
10 Polar Cap~
219 1310 621 0 2 5
0 39 2
0
0 0 1856 0
5 220uF
-16 -18 19 -10
3 C19
-9 -28 12 -20
3 20V
-11 -38 10 -30
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9796 0 0
2
5.89768e-315 5.463e-315
0
7 Ground~
168 1215 675 0 1 3
0 2
0
0 0 53344 0
0
5 GND22
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5952 0 0
2
5.89768e-315 5.46559e-315
0
11 Regulator3~
219 1215 630 0 3 7
0 38 2 39
0
0 0 4928 0
6 KA7810
-21 -28 21 -20
2 U6
-7 -38 7 -30
0
0
14 %D %1 %2 %3 %S
0
0
6 TO-220
7

0 1 2 3 1 2 3 0
88 0 0 0 1 0 0 0
1 U
3649 0 0
2
5.89768e-315 5.46818e-315
0
2 +V
167 1143 585 0 1 3
0 40
0
0 0 53728 0
2 5V
-6 -19 8 -11
2 V7
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3716 0 0
2
42619.7 28
0
7 Ground~
168 1089 756 0 1 3
0 2
0
0 0 53344 0
0
5 GND20
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4797 0 0
2
42619.7 29
0
10 Capacitor~
219 1116 702 0 2 5
0 2 40
0
0 0 832 0
4 10uF
-14 -18 14 -10
3 C18
-11 -28 10 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4681 0 0
2
42619.7 30
0
7 Ground~
168 1341 756 0 1 3
0 2
0
0 0 53344 0
0
5 GND19
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9730 0 0
2
42619.7 31
0
6 IDC40~
219 1231 742 0 40 81
0 22 40 21 40 44 50 20 51 19
52 4 53 3 54 43 55 42 56 18
57 41 58 17 59 60 61 62 63 64
65 66 39 67 2 68 2 69 2 70
2
0
0 0 7776 90
0
2 W2
-113 -13 -99 -5
3 LCD
-117 -3 -96 5
0
0
0
0
5 IDC40
81

0 -9633088 -134323 -9633087 -207977 -9633086 6 -9633085 8 -9633084
10 -9633083 12 -9633082 14 -9633081 16 -211628 18 -781048372
20 -546167348 22 -3177 24 25 26 27 28 29
30 31 -14060019 33 -13588655 35 -195123 37 -195123 39
-195123 -9633088 -134323 -9633087 -207977 -9633086 6 -9633085 8 -9633084
10 -9633083 12 -9633082 14 -9633081 16 -211628 18 -781048372
20 -546167348 22 -3177 24 25 26 27 28 29
30 31 -14060019 33 -13588655 35 -195123 37 -195123 39
-195123 0
0 0 0 512 1 1 0 0
1 J
9874 0 0
2
42619.7 32
0
7 MCP2561
94 744 945 0 8 17
0 37 2 35 36 32 33 34 2
7 MCP2561
1 0 4736 512
7 MCP2561
-25 -37 24 -29
2 U1
-7 -25 7 -17
0
0
0
0
0
4 DIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 0 1 0 0 0
1 U
364 0 0
2
42619.7 33
0
7 MCP2515
94 915 963 0 18 37
0 36 37 71 72 73 74 30 31 2
75 76 77 7 8 9 10 78 35
7 MCP2515
2 0 4736 0
0
2 U7
-3 -43 11 -35
0
0
0
0
0
5 DIP18
37

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 1
2 3 4 5 6 7 8 9 10 11
12 13 14 15 16 17 18 0
0 0 0 512 1 0 0 0
1 U
3656 0 0
2
42619.7 34
0
10 dsPIC33EV~
94 1077 1125 0 28 57
0 6 10 17 22 21 44 20 2 13
14 19 79 5 4 3 43 80 81 2
12 7 8 9 42 18 41 82 11
10 dsPIC33EV~
3 0 4864 512
9 dsPIC33EV
-26 -82 37 -74
2 U4
-3 -70 11 -62
0
0
0
0
0
5 DIP28
57

0 1 2 3 4 5 6 7 8 9
10 11 12 13 14 15 16 17 18 19
20 21 22 23 24 25 26 27 28 1
2 3 4 5 6 7 8 9 10 11
12 13 14 15 16 17 18 19 20 21
22 23 24 25 26 27 28 0
0 0 0 512 1 0 0 0
1 U
3131 0 0
2
42619.7 35
0
9 Resistor~
219 1269 1035 0 2 5
0 6 15
0
0 0 864 0
3 300
-10 -14 11 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 74015272
82 0 0 0 1 0 0 0
1 R
6772 0 0
2
42619.7 36
0
9 Resistor~
219 1323 1035 0 4 5
0 15 5 0 1
0
0 0 864 0
3 10k
-10 -14 11 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 74078176
82 0 0 0 1 0 0 0
1 R
9557 0 0
2
42619.7 37
0
9 Resistor~
219 1615 700 0 3 5
0 26 27 1
0
0 0 864 0
3 220
-10 -12 11 -4
2 R3
-7 -21 7 -13
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5789 0 0
2
5.89768e-315 5.47077e-315
0
110
1 3 2 0 0 4096 0 1 2 0 0 3
1413 1227
1413 1152
1431 1152
0 4 3 0 0 4096 0 0 2 35 0 2
1197 1161
1431 1161
5 0 4 0 0 4096 0 2 0 0 109 2
1431 1170
1188 1170
2 0 5 0 0 4096 0 2 0 0 32 2
1431 1143
1350 1143
0 1 6 0 0 8320 0 0 2 26 0 3
1242 1035
1242 1134
1431 1134
21 13 7 0 0 8320 0 68 67 0 0 4
1044 1134
981 1134
981 981
956 981
14 22 8 0 0 8320 0 67 68 0 0 4
956 972
990 972
990 1125
1044 1125
15 23 9 0 0 8320 0 67 68 0 0 4
956 963
999 963
999 1116
1044 1116
16 2 10 0 0 4224 0 67 68 0 0 4
956 954
1134 954
1134 1080
1118 1080
1 0 2 0 0 0 0 4 0 0 11 2
1260 1206
1260 1215
1 0 2 0 0 8192 0 3 0 0 19 3
1314 1206
1314 1215
1233 1215
2 0 5 0 0 0 0 4 0 0 32 2
1260 1188
1260 1179
2 0 5 0 0 0 0 3 0 0 32 2
1314 1188
1314 1179
1 28 11 0 0 8320 0 5 68 0 0 4
1062 1017
1035 1017
1035 1071
1044 1071
0 2 5 0 0 4224 0 0 5 32 0 4
1350 999
1116 999
1116 1017
1098 1017
1 0 2 0 0 0 0 6 0 0 18 3
972 1179
972 1197
990 1197
20 2 12 0 0 4224 0 68 6 0 0 3
1044 1143
972 1143
972 1161
1 19 2 0 0 0 0 7 68 0 0 3
990 1209
990 1152
1044 1152
1 8 2 0 0 8320 0 8 68 0 0 3
1233 1227
1233 1134
1118 1134
9 0 13 0 0 8320 0 68 0 0 23 5
1118 1143
1170 1143
1170 1233
1188 1233
1188 1269
0 10 14 0 0 4224 0 0 68 22 0 3
1125 1269
1125 1152
1118 1152
1 2 14 0 0 0 0 13 11 0 0 3
1148 1269
1125 1269
1125 1278
2 2 13 0 0 0 0 12 13 0 0 3
1188 1278
1188 1269
1170 1269
1 1 2 0 0 0 0 9 12 0 0 2
1188 1296
1188 1296
1 1 2 0 0 0 0 10 11 0 0 2
1125 1296
1125 1296
1 1 6 0 0 0 0 69 68 0 0 4
1251 1035
1215 1035
1215 1071
1118 1071
2 0 5 0 0 0 0 70 0 0 32 2
1341 1035
1350 1035
1 0 15 0 0 4096 0 15 0 0 29 2
1296 1044
1296 1035
1 2 15 0 0 4224 0 70 69 0 0 2
1305 1035
1287 1035
2 2 16 0 0 4224 0 16 15 0 0 2
1296 1089
1296 1078
1 1 2 0 0 0 0 14 16 0 0 2
1296 1107
1296 1107
13 1 5 0 0 0 0 68 17 0 0 3
1118 1179
1350 1179
1350 972
3 23 17 0 0 16512 0 68 65 0 0 5
1118 1089
1224 1089
1224 954
1242 954
1242 756
25 19 18 0 0 12416 0 68 65 0 0 5
1044 1098
1017 1098
1017 936
1224 936
1224 756
15 13 3 0 0 16512 0 68 65 0 0 5
1044 1188
1035 1188
1035 1215
1197 1215
1197 756
11 9 19 0 0 8320 0 68 65 0 0 3
1118 1161
1179 1161
1179 756
7 7 20 0 0 8320 0 68 65 0 0 3
1118 1125
1170 1125
1170 756
5 3 21 0 0 8320 0 68 65 0 0 3
1118 1107
1152 1107
1152 756
4 1 22 0 0 8320 0 68 65 0 0 3
1118 1098
1143 1098
1143 756
1 0 23 0 0 4224 0 54 0 0 41 2
711 792
711 828
2 2 23 0 0 0 0 20 19 0 0 3
689 828
711 828
711 837
9 1 24 0 0 8320 0 52 20 0 0 3
647 850
666 850
666 828
1 1 2 0 0 0 0 18 19 0 0 2
711 855
711 855
0 2 2 0 0 0 0 0 21 52 0 4
1893 759
1975 759
1975 700
1959 700
1 0 25 0 0 4096 0 21 0 0 51 2
1939 700
1894 700
1 0 26 0 0 4096 0 71 0 0 60 2
1597 700
1585 700
2 0 2 0 0 0 0 22 0 0 61 4
1654 700
1669 700
1669 760
1584 760
1 2 27 0 0 4224 0 22 71 0 0 2
1634 700
1633 700
1 0 25 0 0 0 0 24 0 0 51 2
1840 727
1840 718
2 0 25 0 0 0 0 25 0 0 51 2
1894 727
1894 718
3 1 25 0 0 4224 0 30 23 0 0 3
1823 718
1894 718
1894 691
0 1 2 0 0 0 0 0 25 53 0 3
1840 759
1894 759
1894 745
2 0 2 0 0 0 0 24 0 0 56 3
1840 744
1840 759
1795 759
0 2 28 0 0 4096 0 0 26 57 0 2
1741 718
1741 727
1 1 2 0 0 0 0 28 26 0 0 2
1741 766
1741 745
1 2 2 0 0 0 0 27 30 0 0 2
1795 766
1795 751
1 1 28 0 0 4224 0 29 30 0 0 3
1741 691
1741 718
1767 718
1 0 26 0 0 0 0 37 0 0 60 2
1531 728
1531 719
2 0 26 0 0 0 0 36 0 0 60 2
1585 728
1585 719
3 1 26 0 0 4224 0 31 38 0 0 3
1514 719
1585 719
1585 692
0 1 2 0 0 0 0 0 36 62 0 3
1531 760
1585 760
1585 746
2 0 2 0 0 0 0 37 0 0 65 3
1531 745
1531 760
1486 760
0 2 29 0 0 4096 0 0 35 66 0 2
1432 719
1432 728
1 1 2 0 0 0 0 33 35 0 0 2
1432 767
1432 746
1 2 2 0 0 0 0 34 31 0 0 2
1486 767
1486 752
1 1 29 0 0 4224 0 32 31 0 0 3
1432 692
1432 719
1458 719
1 1 2 0 0 0 0 40 41 0 0 2
810 1089
810 1089
1 1 2 0 0 0 0 39 42 0 0 2
873 1089
873 1089
0 7 30 0 0 8320 0 0 67 72 0 3
810 1053
810 990
882 990
0 8 31 0 0 4224 0 0 67 71 0 3
873 1053
873 999
882 999
2 2 31 0 0 0 0 42 43 0 0 3
873 1071
873 1053
855 1053
2 1 30 0 0 0 0 41 43 0 0 3
810 1071
810 1053
833 1053
1 2 2 0 0 0 0 44 45 0 0 2
684 1017
684 1010
1 5 32 0 0 4224 0 45 66 0 0 3
684 990
684 963
711 963
8 0 2 0 0 0 0 66 0 0 86 4
711 936
702 936
702 981
783 981
6 6 33 0 0 8320 0 52 66 0 0 4
647 877
684 877
684 954
711 954
7 7 34 0 0 8320 0 66 52 0 0 4
711 945
693 945
693 868
647 868
2 0 35 0 0 4096 0 47 0 0 80 2
864 891
864 882
1 1 2 0 0 0 0 46 47 0 0 2
864 909
864 909
0 18 35 0 0 4224 0 0 67 83 0 4
801 882
972 882
972 936
956 936
2 0 35 0 0 0 0 49 0 0 83 3
747 873
747 864
801 864
1 1 2 0 0 0 0 48 49 0 0 2
747 891
747 891
1 3 35 0 0 0 0 50 66 0 0 3
801 856
801 954
777 954
4 1 36 0 0 12416 0 66 67 0 0 4
777 963
828 963
828 936
882 936
9 0 2 0 0 0 0 67 0 0 86 2
882 1008
783 1008
1 2 2 0 0 0 0 51 66 0 0 3
783 1017
783 945
777 945
1 2 37 0 0 12416 0 66 67 0 0 4
777 936
819 936
819 945
882 945
1 8 2 0 0 0 0 53 52 0 0 3
666 912
666 859
647 859
2 0 38 0 0 4096 0 55 0 0 91 2
1179 630
1179 621
0 1 2 0 0 0 0 0 55 92 0 3
1215 661
1179 661
1179 648
1 1 38 0 0 4224 0 56 60 0 0 3
1179 594
1179 621
1187 621
1 2 2 0 0 0 0 59 60 0 0 2
1215 669
1215 654
1 0 2 0 0 0 0 57 0 0 94 2
1317 666
1341 666
2 0 2 0 0 0 0 58 0 0 107 3
1316 621
1341 621
1341 702
1 0 39 0 0 4096 0 58 0 0 97 2
1299 621
1277 621
2 0 39 0 0 0 0 57 0 0 97 2
1299 666
1278 666
3 32 39 0 0 8320 0 60 65 0 0 3
1243 621
1278 621
1278 721
34 0 2 0 0 0 0 65 0 0 99 3
1287 721
1287 702
1296 702
36 0 2 0 0 0 0 65 0 0 101 3
1296 721
1296 702
1305 702
4 0 40 0 0 4096 0 65 0 0 104 3
1152 721
1152 675
1143 675
38 0 2 0 0 0 0 65 0 0 107 3
1305 721
1305 702
1314 702
21 26 41 0 0 8320 0 65 68 0 0 5
1233 756
1233 945
1026 945
1026 1089
1044 1089
17 24 42 0 0 8320 0 65 68 0 0 5
1215 756
1215 927
1008 927
1008 1107
1044 1107
1 0 40 0 0 4224 0 61 0 0 105 2
1143 594
1143 702
2 2 40 0 0 0 0 63 65 0 0 3
1125 702
1143 702
1143 721
1 1 2 0 0 0 0 63 62 0 0 3
1107 702
1089 702
1089 750
1 40 2 0 0 0 0 64 65 0 0 4
1341 750
1341 702
1314 702
1314 720
15 16 43 0 0 4224 0 65 68 0 0 5
1206 756
1206 1224
1026 1224
1026 1179
1044 1179
11 14 4 0 0 4224 0 65 68 0 0 3
1188 756
1188 1188
1118 1188
5 6 44 0 0 4224 0 65 68 0 0 3
1161 756
1161 1116
1118 1116
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
